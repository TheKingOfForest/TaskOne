`timescale 1ns/1ps
module alu_test;

reg[31:0] instruction, regA, regB;
wire[31:0] result;
wire[2:0] flag;

alu testalu(instruction, regA, regB, result, flag);

initial begin
    $dumpfile("test_ALU.vcd");
    $dumpvars(0,instruction, regA, regB, result, flag);
end

initial begin
    $display("instruction|regA|regB|result|flag");
    $monitor("%b  %b  %b  %b  %b",instruction, regA, regB, result, flag);
    #10 $display("-----------+--+----+----+--------+--add---+--------+-----+--------+--------");
            // 1 + 2 = 3 general
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // negtive test
            // -2 + 1 = -1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;
            // overflow flag test (positive)
            // 32'h7FFFF_FFFF + 32'd1 = 32'hFFFF_FFFF
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
            regA <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // overflow flag test (negative)
            // 32'h8000_0000 + 32'hFFFF_FFFF = 33'h1_7FFF_FFFF
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
            regA <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
            regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
        #10 $display("-----------+--+----+----+--------+--addi--+--------+-----+--------+--------");
            // 1 + 8 = 9 general
            #10 instruction <= 32'b0010_0000_0000_0000_0000_0000_0000_1000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // negtive test
            // -2 + 1 = -1
            #10 instruction <= 32'b0010_0000_0000_0000_0000_0000_0000_0001;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;
            // negative imme test
            // -1 + 2 = 1
            #10 instruction <= 32'b0010_0000_0000_0000_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // overflow flag test (positive)
            // 32'h7FFFF_FFFF + 32'd1 = 32'hFFFF_FFFF
            #10 instruction <= 32'b0010_0000_0000_0000_0000_0000_0000_0001;
            regA <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
            // overflow flag test (negative)
            // 32'h8000_0000 + 32'hFFFF_FFFF = 33'h1_7FFF_FFFF
            #10 instruction <= 32'b0010_0000_0000_0000_1111_1111_1111_1111;
            regA <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        #10 $display("-----------+--+----+----+--------+--addu--+--------+-----+--------+--------");
            // 1 + 2 = 3
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0001;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        #10 $display("-----------+--+----+----+--------+--addiu-+--------+-----+--------+--------");
            // 1 + 15 = 16
            #10 instruction <= 32'b0010_0100_0000_0000_0000_0000_0000_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // unsigned extension test
            // 65535 + 1 = 65536
            #10 instruction <= 32'b0010_0100_0000_0000_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--sub---+--------+-----+--------+--------");
            // 2 - 1 = 1 general
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // (-1) - (-2) = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
            regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;
            // negative test
            // 0 - 1 = -1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // overflow flag test
            // 32'h7FFF_FFF - (-1) = 32'h8000_0000
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
            regA <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
            regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
            // overflow flag test
            // 32'h8000_000 - 1 = 33'h1_7FFF_FFFF
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
            regA <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--subu--+--------+-----+--------+--------");
            // 2 - 1 = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // zero flag test
            // 1 - 1 = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--and---+--------+-----+--------+--------");
            // 3 & 5 = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0100;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        #10 $display("-----------+--+----+----+--------+--andi--+--------+-----+--------+--------");
            // 3 & 5 = 1
            #10 instruction <= 32'b0011_0000_0000_0001_0000_0000_0000_0011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
            // unsigned externsion test
            // 32'hFFFF_FFFF & 65535 = 65535
            #10 instruction <= 32'b0011_0000_0000_0001_1111_1111_1111_1111;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
        #10 $display("-----------+--+----+----+--------+--nor---+--------+-----+--------+--------");
            // ~(3 | 5) = 32'hFFFF_FFF8
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        #10 $display("-----------+--+----+----+--------+--or----+--------+-----+--------+--------");
            // 3 | 5 = 7
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0101;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        #10 $display("-----------+--+----+----+--------+--ori---+--------+-----+--------+--------");
            // 3 | 5 = 7
            #10 instruction <= 32'b0011_0100_0000_0001_0000_0000_0000_0011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
            // unsigned externsion test
            // 0 & 65535 = 65535
            #10 instruction <= 32'b0011_0100_0000_0001_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        #10 $display("-----------+--+----+----+--------+--xor---+--------+-----+--------+--------");
            // 3 ^ 5 = 6
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_0110;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        #10 $display("-----------+--+----+----+--------+--xori--+--------+-----+--------+--------");
            // 3 ^ 5 = 6
            #10 instruction <= 32'b0011_1000_0000_0001_0000_0000_0000_0011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;
            // unsigned externsion test
            // 32'h0000_0000 & 65535 = 65535
            #10 instruction <= 32'b0011_1000_0000_0001_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        #10 $display("-----------+--+----+----+--------+--beq---+--------+-----+--------+--------");
            // equal test
            #10 instruction <= 32'b0001_0000_0000_0001_0000_0000_0000_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // inequal test
            #10 instruction <= 32'b0001_0000_0000_0001_0000_0000_0000_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--bne---+--------+-----+--------+--------");
            // equal test
            #10 instruction <= 32'b0001_0100_0000_0001_0000_0000_0000_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // inequal test
            #10 instruction <= 32'b0001_0100_0000_0001_0000_0000_0000_0000;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--slt---+--------+-----+--------+--------");
            // 1 < 2
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // 2 > 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // 1 = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // slt test (signed test)
            // -1 < 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1010;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--slti--+--------+-----+--------+--------");
            // 1 < 2
            #10 instruction <= 32'b0010_1000_0000_0000_0000_0000_0000_0010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001; 
            // 2 > 1
            #10 instruction <= 32'b0010_1000_0000_0000_0000_0000_0000_0001;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // 1 = 1
            #10 instruction <= 32'b0010_1000_0000_0000_0000_0000_0000_0001;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // slti test (signed test)
            // 1 > -1
            #10 instruction <= 32'b0010_1000_0000_0000_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--sltu--+--------+-----+--------+--------");
            // 1 < 2
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // 2 > 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // sltu test - 0 
            // 1 = 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // sltu test (unsigned test)
            // 32'hFFFF_FFFF > 1
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
            regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // sltu test (unsigned test)
            // 1 < 32'hFFFF_FFFF
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
        #10 $display("-----------+--+----+----+--------+--sltiu-+--------+-----+--------+--------");
        // sltiu rt, rs, imm - 0xb, rs, rt, imm
            // sltiu test - 1 (negative flag)
            // 1 < 2
            #10 instruction <= 32'b0010_1100_0000_0000_0000_0000_0000_0010;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // sltiu test - 0 
            // 2 > 1
            #10 instruction <= 32'b0010_1100_0000_0000_0000_0000_0000_0001;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            // sltiu test (zero flag)
            // 1 = 1
            #10 instruction <= 32'b0010_1100_0000_0000_0000_0000_0000_0001;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            // sltu test (unsigned test)
            // 32'hFFFF_FFFF > 1
            #10 instruction <= 32'b0010_1100_0000_0000_0000_0000_0000_0001;
            regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
            // sltu test (unsigned test)
            // 1 < 32'h0000_FFFF
            #10 instruction <= 32'b0010_1100_0000_0000_1111_1111_1111_1111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        #10 $display("-----------+--+----+----+--------+--lw----+--------+-----+--------+--------");
        // lw rt, rs(offset) - 0x23, rs, rt, offset
            // lw test
            // 32'h0008_0000 + 80
            #10 instruction <= 32'b1000_1100_0000_0000_0000_0000_0101_0000;
            regA <= 32'b0000_0000_0000_1000_0000_0000_0000_0000;
            // 32'h0008_0000 - 80 (signed extension)
            #10 instruction <= 32'b1000_1100_0000_0000_1111_1111_1011_0000;
            regA <= 32'b0000_0000_0000_1000_0000_0000_0000_0000;
        #10 $display("-----------+--+----+----+--------+--sw----+--------+-----+--------+--------");
        // sw rt, rs(offset) - 0x2b, rs, rt, offset
            // sw test
            // 32'h0008_0000 + 80
            #10 instruction <= 32'b1010_1100_0000_0000_0000_0000_0101_0000;
            regA <= 32'b0000_0000_0000_1000_0000_0000_0000_0000;
            // 32'h0008_0000 - 80 (signed extension)
            #10 instruction <= 32'b1010_1100_0000_0000_1111_1111_1011_0000;
            regA <= 32'b0000_0000_0000_1000_0000_0000_0000_0000;
        #10 $display("-----------+--+----+----+--------+--sll---+--------+-----+--------+--------");
            // 32'h1234_5678 << 4 = 32'h2345_6780
            #10 instruction <= 32'b0000_0000_0000_0000_0000_0001_0000_0000;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
        #10 $display("-----------+--+----+----+--------+--sllv--+--------+-----+--------+--------");
            // 32'h1234_5678 << 4 = 32'h2345_6780
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0100;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
            // the least five bits test
            // 32'h1234_5678 << 4 = 32'h2345_6780
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0100;
            regA <= 32'b1111_1111_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
        #10 $display("------------------------------------srl---+--------+-----+--------+--------");
            // 32'h1234_5678 >> 4 = 32'h0123_4567
            #10 instruction <= 32'b0000_0000_0000_0000_0000_0001_0000_0010;
            regA <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
        #10 $display("-----------+--+----+----+--------+--srlv--+--------+-----+--------+--------");
            // 32'h1234_5678 >> 4 = 32'h0123_4567
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0110;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
            // the least five bits test
            // 32'h1234_5678 >> 4 = 32'h0123_4567
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0110;
            regA <= 32'b1111_1111_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
        #10 $display("-----------+--+----+----+--------+--sra---+--------+-----+--------+--------");
            // 32'h1234_5678 >>> 4 = 32'h023_4567
            #10 instruction <= 32'b0000_0000_0000_0000_0000_0001_0000_0011;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
            // 32'h8765_4321 >>> 4 = 32'hF876_5432 (negative flag)
            #10 instruction <= 32'b0000_0000_0000_0000_0000_0001_0000_0011;
            regB <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
        #10 $display("-----------+--+----+----+--------+--srav--+--------+-----+--------+--------");
            // 32'h1234_5678 >>> 4 = 32'h0123_4567
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
            // 32'h8765_4321 >>> 4 = 32'F876_5432
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0111;
            regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            regB <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
            // the least five bits
            // 32'h1234_5678 >>> 4 = 32'h0123_4567
            #10 instruction <= 32'b0000_0000_0000_0001_0000_0000_0000_0111;
            regA <= 32'b1111_0000_0000_0000_0000_0000_0000_0100;
            regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;
    #10 $finish;
end

endmodule